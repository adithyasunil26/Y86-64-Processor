module decode(

)
  
endmodule