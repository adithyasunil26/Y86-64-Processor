module fetch(
  clk,
)

endmodule