module decode(
  
)

endmodule