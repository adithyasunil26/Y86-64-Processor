`timescale 1ns / 1ps

module decode(

)



endmodule