`timescale 1ns / 1ps

module and1x1(
  input a,
  input b,
  output ans
  );

  and g1(ans,a,b);
  
endmodule