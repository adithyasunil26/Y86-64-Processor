module fetch(

)

endmodule