`timescale 1ns / 1ps

module not1x1(
  input a,
  output ans
  );

  not g1(ans,a);  

endmodule